`ifndef ALU_DEFS_SVH
`define ALU_DEFS_SVH

/*
    This header defines common data structrue & constants in alu module
*/

// nmc defs
`include "nmc_defs.svh"

`endif
