// alveo_cim
`include "common_defs.svh"

module alveo_cim #(

) (

);

// TODO

endmodule
