`ifndef COMMON_DEFS_SVH
`define COMMON_DEFS_SVH

/*
    This header defines common data structrue & constants in the whole soc
*/

// project configuration
`default_nettype wire
`timescale 1ns / 1ps

// compile_options
`include "compile_options.svh"

`endif
