`ifndef ALU_DEFS_SVH
`define ALU_DEFS_SVH

/*
    This header defines common data structrue & constants in alu module
*/

// cim defs
`include "cim_defs.svh"

`endif
