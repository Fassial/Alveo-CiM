`ifndef CAM_DEFS_SVH
`define CAM_DEFS_SVH

/*
    This header defines common data structrue & constants in cam module
*/

// common defs
`include "common_defs.svh"

`endif
