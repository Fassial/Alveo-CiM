`ifndef CIM_DEFS_SVH
`define CIM_DEFS_SVH

/*
    This header defines common data structrue & constants in cim module
*/

// common defs
`include "common_defs.svh"

`endif
